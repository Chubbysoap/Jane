`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/17/2025 08:54:59 AM
// Design Name: 
// Module Name: tb_parse_vectors
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// SystemVerilog Testbench for Parsing "R10 L798" into Vectors
module tb_parse_vectors;

    // Declare vectors as unpacked arrays
    logic [0:0] direction [1:0];  // 1-bit per direction (0 or 1)
    logic [31:0] magnitude [1:0]; // 32-bit for magnitudes (adjust if needed)

    initial begin
        // Input string
        string input_str = "R41 R17 L15 L2 L41 L47 L42 R8 R29 L32 L14 R26 R28 L35 R2 L4
L27
R37
L14
R2
R50
R12
L13
L3
L29
L37
L6
R43
R13
L26
L24
R23
R29
R18
R8
R20
R50
L23
L24
R25
R31
R6
L19
L25
R6
L43
R21
L15
R3
L38
R94
L11
R27
R38
R19
L73
L94
L9
R74
R73
L23
R93
R92
R40
R17
L57
L33
R53
L98
L25
L71
L26
R89
L30
R66
L88
L37
L42
L58
L53
L40
L7
R96
L56
R60
L59
L14
L11
L49
L24
R38
R19
L62
L38
L93
L7
R30
R31
L3
L13
R9
L563
R75
R34
L4
L34
L162
L3
R146
L97
R94
L49
L99
L992
R93
R4
L6
L91
L27
R86
R50
R66
R57
L59
R27
L38
R15
R23
L65
L77
L996
R98
L6
R27
L929
R103
L78
L77
R80
R972
L94
L36
R7
R28
R43
L72
R72
L621
L323
L56
R87
R23
L110
L93
L731
R42
L18
L9
R9
L72
R9
R14
R69
R34
L454
L41
L82
R7
L66
R5
L672
R31
L13
R531
R89
R31
L25
L73
L922
L47
L316
R13
R84
L34
R647
R92
L8
R69
R135
R60
R5
L464
L99
R63
L19
R907
L78
R90
R38
R62
R66
L466
R462
L762
L287
R678
L91
R72
R81
L356
L859
R63
L28
L69
L4
L877
L23
L1
L2
L897
L54
L49
R15
R89
R10
L21
R11
L46
L832
R57
L43
L70
L859
L8
R19
R81
L32
R1
L83
R33
L19
R19
L19
R10
L27
L83
L57
L57
R14
R31
L97
R66
R147
L747
L52
R392
L65
R97
L99
R20
R13
L80
L43
L90
L190
R797
L89
R992
R997
L89
L37
R77
R49
R86
R214
L13
L689
R17
R59
L48
L24
R98
L74
R15
L766
L670
L5
R645
L445
L76
R76
R53
L60
L93
R71
R668
L39
R450
R288
R76
L14
R9
L9
R43
L66
R67
R572
L63
R658
R89
L18
R747
L211
R13
R41
L44
L16
R188
L576
R76
L464
R364
L154
L38
R65
R2
L70
L705
L56
R256
L56
L44
L5
L95
L897
L16
L19
L647
R4
L78
L80
R58
L75
L50
R16
R614
R70
L48
R48
L47
R74
L38
L89
R548
R52
R23
L22
L20
R274
R525
L82
L76
L90
R68
L649
L61
R12
L97
R95
L10
R510
R274
R26
L34
L66
R18
L25
L54
R29
R32
R59
R578
L937
R91
L252
R84
R77
R27
R77
L26
R3
L81
R91
L40
L23
L81
R753
L78
L338
R9
R1
R873
R10
R85
R80
R358
R45
R430
L3
L60
R621
R67
R69
R56
R97
L51
R183
L580
R69
L79
R68
R811
R57
R7
L14
L29
R36
L391
L109
L2
R2
L95
R18
L23
L79
R79
L71
R696
L34
R73
R528
L782
R271
R29
L310
L17
L383
R59
R75
R84
R162
R520
R92
R266
R363
R247
L32
L50
L86
L27
L73
L7
R880
R331
R96
L35
L65
R42
R34
L176
L372
L54
R26
L64
R64
R412
R83
L95
R22
R78
R60
R54
L14
R85
L985
L57
R72
L15
L2
R51
L24
R38
L3
R93
L53
R73
R16
R44
L33
L46
L305
R51
L77
L18
L795
R361
L64
R353
L88
L598
R6
L50
L24
R94
R87
L916
L45
L26
L630
L18
L52
L75
R7
L32
R25
R75
L75
R35
L60
L70
R70
R34
R36
L87
R94
R23
L67
R667
R16
R84
L8
R96
L26
R84
R54
L61
L15
L48
R63
L49
L10
R37
R183
R951
L51
L342
R208
R695
L61
R80
R20
L80
L570
L350
R40
L922
R703
L61
R40
R760
R703
R40
L3
L842
R976
L53
R98
R49
L75
R64
L17
R89
R65
L54
R2
R98
R896
L96
R49
R651
L15
R15
R64
R14
L78
R86
R3
R39
R172
L69
R70
L601
R18
L307
L11
L59
L41
L92
L8
R78
R107
L85
L90
L10
L6
L994
R27
R30
R43
L139
L7
R46
L2
R2
L719
R58
L39
L948
L52
R29
L91
L46
L92
R42
L58
L84
L31
L29
L65
R41
L110
L81
L64
L50
L74
L98
R61
R73
L73
L3
L621
L876
R25
L49
R8
R16
L58
L91
L988
R37
L82
R82
L55
R558
L22
L90
L91
R94
R6
L92
L8
L99
L1
R97
R105
R741
L70
R94
L85
R577
R11
R730
L291
L9
R48
R1
L630
L10
R85
R218
L12
L347
L53
R664
L57
L65
L42
L90
L93
L859
R48
R394
R60
L49
R63
L55
R20
L5
R17
R19
R30
L75
L21
L50
L40
R86
R15
R22
R983
R12
L32
R4
L4
L48
L16
L83
L25
L49
L86
L93
L34
L40
R185
L11
R54
L29
L826
L75
R1
L47
R122
L64
L36
L22
R59
L80
L257
L80
R1
L621
R25
L84
R2
R57
R61
R39
R474
R26
R291
L50
R15
R39
R2
L56
L41
R695
L160
R95
R46
L76
L95
R95
R9
R361
R3
R722
R86
L81
L73
L87
L553
R66
L71
R934
L60
R37
L59
R75
R54
L692
R45
R84
R23
L12
R66
R23
R925
L66
R46
R7
R88
R32
L97
L19
R35
R45
L96
R53
L454
L98
L101
L85
R85
L20
L646
L94
R370
L10
L90
L45
R940
R95
R15
R561
R80
R44
L25
R89
L64
L20
L893
L87
R65
L32
R42
R25
L328
L76
L79
L17
R327
L27
L27
L551
R12
R881
L71
L96
R89
R63
L57
L94
R93
L42
L54
L31
R483
R102
R89
R59
R24
L60
L12
R62
R38
L21
R21
R74
R20
R6
R20
R72
L37
L55
L63
L37
R96
R63
L59
L14
R82
L468
L51
R25
R26
R44
R57
L72
R923
R80
R99
L66
L265
L94
L73
R466
L99
L27
R27
R30
L67
R33
R31
R88
R255
L70
R627
R383
R724
R99
L911
R53
R81
R19
R94
L983
L56
R70
L87
L85
R31
L23
R464
L63
L63
R26
L65
L37
L98
L234
L66
L378
R122
L64
R20
L31
R822
R9
L68
R68
R74
L42
R928
R979
R61
R678
L78
R75
L475
L85
R7
L31
L91
L62
L85
R71
L84
L35
L34
R40
L11
R88
R87
R42
R57
L58
L716
R34
R60
R206
L38
R72
L39
L20
L95
L234
R476
R57
R221
R44
L44
R522
R49
L71
R13
L495
R20
L83
R45
R81
L56
L25
R14
R976
R340
R82
L12
L34
L77
R460
L38
R86
L97
L60
L530
R80
R49
L39
R74
R847
L7
L57
R52
R86
R8
L3
R37
L37
L58
L42
L947
R47
L5
R805
R47
R53
L81
R4
L93
R91
R70
L91
L15
L485
R15
L15
L42
R4
L50
R473
L66
R99
L96
R4
L26
R58
R3
L78
R38
L8
R61
R21
L48
L47
R34
R20
R81
L32
L3
L40
R93
R79
L70
R15
L72
L99
L71
R25
R40
L19
L78
L3
R79
R19
R11
R691
R619
R81
L95
L55
R41
R9
R636
L75
L7
L94
R740
R64
R36
R32
R68
R332
R68
R14
R81
L12
R11
R6
L38
R70
L397
R68
L47
L87
R31
L75
R49
R87
L13
L92
R46
L602
R58
L58
R692
L456
R98
L92
R58
R65
L565
R49
L73
L763
R660
R96
L17
R16
R74
L542
L19
L20
L48
L13
L28
R28
L18
R52
R66
R61
L94
R33
R55
L55
L45
R70
L51
R26
R383
R17
L96
R28
R98
L20
R875
L77
L208
R27
L128
L199
L38
R43
L38
L69
R28
L24
L17
R99
L84
R42
L95
L56
L148
L66
R4
R16
L95
L261
R18
R53
L12
L628
L72
L81
R59
L36
R46
L23
L65
R12
R2
L79
R65
R89
R34
R8
L31
L12
L5
R77
L37
L46
L426
R49
L41
L37
L36
L86
L667
L82
R88
R764
L3
R333
L7
L40
L86
R679
R796
L29
L46
R737
L37
R53
L89
L64
R63
L63
L38
R838
L58
L42
L55
R55
L64
R99
R72
L392
L75
R560
R88
L64
R76
R77
L82
L61
L94
R82
L76
L96
L273
L29
R18
L66
R74
L877
R73
R52
L22
R21
L80
L59
L23
L430
L429
L73
R73
L1
L995
L638
R419
L71
R75
R10
R601
R63
L63
R98
L32
L21
R55
R37
L535
R98
L75
R722
R89
L36
R90
R7
L35
L62
R34
R62
L32
L18
L46
R880
L84
R4
L81
R44
R86
L49
L131
L69
R587
L87
L65
R18
R64
R98
R884
R50
R14
R8
R29
L71
R54
L21
L362
R49
L57
L79
R74
R13
R280
L597
R17
R67
R37
R96
L35
L83
L82
L28
R28
L48
R48
L91
R70
R68
L47
L54
L21
L25
L137
L49
R20
R66
L95
L5
R86
R89
R61
R910
L46
R90
L60
L84
L16
L28
L362
L940
L75
R93
L820
L99
L9
L93
R45
R34
R324
R94
L194
L77
R77
R34
L34
R89
R267
L45
L15
L89
R79
R52
R74
R88
R18
L57
R89
L50
R89
R58
L85
L45
R71
R12
R344
R51
R17
L14
R25
R62
R12
R703
R38
R362
L90
L10
L656
L735
R57
R94
L60
L90
L49
L33
R92
L77
L43
R91
L51
R62
L2
L34
L25
R28
R31
R8
R44
R86
L224
L78
R64
R89
L89
L55
R99
L28
L20
L33
L63
L60
L562
L21
L557
L87
L84
R9
R81
L696
R91
R95
R91
L26
L74
R15
L15
L60
L40
R8
R92
L89
L76
L67
L468
L360
R65
L5
R80
L80
L33
R98
R31
R104
L32
R152
L17
L3
R1
L337
R67
L33
R83
R719
L30
R189
R34
L93
R31
R669
R28
L56
R28
R55
R45
L93
L7
R72
R29
L951
L1
L31
R615
R18
L17
L23
R89
R70
R47
R83
L18
R18
R4
L4
R88
R77
L65
R54
R51
R33
R74
R65
R30
L15
R94
L186
L912
L95
R477
R87
L257
R24
R22
L46
R70
L70
R58
L682
R24
L58
R40
R18
R6
L6
L62
R34
R75
R53
L628
L179
R7
L92
R92
L21
R53
L63
L50
L219
L4
R14
R90
R53
R15
L68
R18
R82
L82
R91
R91
L41
R41
L923
R23
L98
L15
R67
R81
R24
L40
L19
L689
R8
R17
R38
L66
L8
R73
R30
R35
R909
L447
L72
R72
L527
R7
R27
R78
L86
L99
L65
R79
L45
L61
R93
L223
R36
R77
L91
L81
L419
L37
R72
L35
L63
R31
R96
L44
L20
L219
L84
L69
L34
R79
L74
L34
R35
L12
L88
L38
R838
L882
L919
R22
L680
L41
L88
L85
R23
L50
R57
L57
R77
R99
L976
R60
R40
L72
L28
L17
L16
R78
R49
L30
R136
L735
L65
L39
L961
R16
R83
R73
R18
L90
L36
R36
R552
R48
L937
R37
R37
R4
R233
R26
L70
L30
L98
L2
R8
R44
L52
R14
L663
R49
R93
R907
L36
R36
R589
L11
R1
R927
R98
L4
R35
L435
L6
R817
R3
L314
L41
R941
R61
L34
R795
R62
R382
R46
L87
L25
L91
L63
R54
R10
R88
R669
R733
L7
L93
R43
R97
R1
L77
L64
R12
L331
L581
L13
R13
L21
L79
R17
R42
R41
R3
R97
L977
L923
R54
R30
R16
R82
R71
L53
L821
L46
R567
L386
L287
L54
L56
L17
R93
R98
L91
R8
L8
L20
R20
R88
R48
L475
L158
L90
L15
L75
R37
L260
L44
L44
L584
L34
R98
L92
L67
R50
R26
L11
R2
R180
R80
L578
L13
R31
R72
R52
L9
L91
L94
L30
L82
R86
R196
L326
R92
L66
R24
L24
R30
R170
L13
L96
R9
R2
R998
L9
R47
L57
R319
R13
R29
L2
R18
L658
L25
L35
L10
L79
R71
L22
R641
L20
R16
L57
L80
L391
R91
L12
R712
L64
R811
R53
L95
L66
R90
R78
L7
L45
L55
L102
R2
L454
L31
R1
R98
R86
L76
L28
L54
L86
R16
R128
L972
R472
R19
R81
L41
L687
L34
L91
L183
L364
R42
R8
R508
L10
R20
R743
L53
L12
R854
R35
L35
R578
R538
L16
R37
R71
L8
L79
R79
R77
R723
R66
R34
L6
L40
L54
R24
R24
R43
L76
L72
R57
R59
L85
R49
L32
R39
R48
L78
L99
L98
L99
R96
R11
L94
L45
R85
R843
L819
R19
L88
R88
L20
R417
R3
R51
R49
R69
L69
L4
L412
L46
L5
R38
L44
L63
R265
R37
L67
L84
L33
L104
R302
R64
L16
R72
R80
R461
R83
R76
L4
R83
L34
R966
R615
L35
R248
L441
R903
R42
R46
L14
R25
R708
L47
L61
L602
L72
R29
R88
R27
L761
L227
R705
R13
L85
R180
R8
R97
L97
R38
R59
R11
R606
L48
R9
R305
R17
R66
L16
R13
L63
R9
L47
R38
L363
L37
R11
R88
R98
R3
L33
R88
L555
R80
R17
L97
L453
R28
R256
R92
L23
L42
L51
R854
R39
L8
R67
L52
R704
R84
R518
R66
L18
R13
R26
R70
R30
L371
R16
L98
R36
R989
R16
R59
L747
R12
R53
L245
L143
L77
R67
R193
R40
L53
R53
L24
L452
R3
L22
L45
L60
R82
R18
R14
L79
L17
R9
R26
R47
L247
L781
L72
L9
L85
R23
R534
L63
L808
R20
L46
L250
L316
L708
R8
L70
L42
L1
R62
L263
R11
L84
R87
R38
R210
R52
R28
R72
R81
R19
L34
R88
L402
L452
R2
L64
R65
R19
R78
R5
L11
L49
R55
R10
L14
L96
L69
L2
R88
L58
R41
L79
L21
R89
L97
R708
L207
R61
L54
L68
L27
L85
L2
R18
R60
R4
R812
L84
L15
L13
R78
L31
L12
R46
L42
L14
L51
R66
L40
L411
R11
L46
R978
L91
R59
R19
R38
L57
R1
R99
R70
L899
R48
R53
R3
R82
R459
R8
L80
R58
L2
L60
R360
L43
R743
R97
R833
R72
L84
R88
R63
R10
L33
R2
L21
R6
L328
L18
R331
R81
R60
R82
L36
L78
L55
L40
L21
L78
L18
L15
R82
L122
L63
R3
R3
R89
L92
R456
R44
R11
R54
L8
R43
L574
L10
R84
L28
R685
L62
R905
R50
R91
R59
L36
R354
R82
L226
R9
L83
L80
R290
R34
L721
L47
L76
R451
R49
R51
R81
R34
L366
R33
L50
R17
R52
L49
L3
L426
L63
L65
L946
R92
R37
L29
R75
L475
R1
R67
R61
R86
L37
R34
L39
L27
R254
R414
L29
L52
R96
L829
L74
R56
R34
L65
R329
R55
L59
L43
R67
R52
L653
L43
L56
R73
R37
R6
R80
R504
R63
L759
L30
L65
R58
R33
R304
R20
R85
L14
L10
L658
L6
R79
R78
R22
R75
L159
R35
L791
R669
R571
L25
L62
L13
L39
R112
R73
R54
R549
R39
L83
L45
L75
L19
R661
R37
R14
R22
R10
R90
L909
L863
L28
R36
R8
R811
R45
L81
L19
L92
R92
L868
L732
L47
L5
L48
L31
L89
L80
R642
L986
L41
R217
R11
R69
R88
R979
L79
R37
R48
R15
L33
L67
R14
R60
L87
R19
L6
R981
L81
L33
L71
R13
L719
R36
L31
L95
L94
R23
L88
L41
R17
R73
L90
L29
R89
R84
L59
R7
L66
R41
R71
R62
L50
L76
L618
R44
R78
L44
R66
L61
L39
L64
L98
R62
R440
L78
R38
L48
L50
R683
L40
L21
R76
R71
L71
L63
L53
R84
R332
R94
L8
L32
L44
R90
R7
R93
L637
L821
L87
L17
L83
L6
R51
R4
L74
R70
R185
L36
L208
L41
L16
L34
L85
R28
R7
R903
L3
R289
R11
L98
L2
R1
R99
R88
R12
L34
R96
R12
L74
R23
L23
R44
R54
L19
R21
L25
R804
L10
L13
R44
R67
R738
R56
L43
L18
L25
L47
L28
R13
R954
R733
R80
L35
R55
L56
L26
R682
R5
L73
L71
L61
R57
R724
R35
L3
L54
R741
L27
R84
R43
R689
L89
L31
R23
L8
L84
L55
L45
R34
R66
L995
R26
L7
L50
L640
R66
R92
R55
R4
R835
L36
L14
R201
L5
L58
L265
L31
R22
R6
R94
L90
R69
L79
L29
L831
L404
L70
R94
L60
L367
L426
R693
L429
R305
L20
L56
R56
R44
L49
R649
R15
R985
R277
R923
L56
R902
L24
R412
L34
R27
L75
R48
L98
R98
L65
L35
R39
L39
R19
R445
L54
R90
L81
R81
L52
R52
L32
L814
L15
R38
R21
R35
R28
R39
R97
L781
L10
L53
L53
R385
R758
R1
L35
L35
L74
R32
R73
R11
L79
L437
R13
L46
L87
L80
R13
L39
L774
R64
R306
R30
L61
R661
R166
R34
L122
L78
R63
R33
L96
L51
R51
R65
R26
L63
L906
R778
L726
R73
R53
L63
R784
R83
L4
L26
L56
L9
L99
R80
L90
R677
L77
L13
R13
R33
R267
R98
R52
R250
L59
L44
L97
L86
L72
L42
L454
R54
R4
L15
R42
L42
R10
R1
R28
L88
L16
R76
L28
L75
L97
R45
R55
L29
R29
R18
R55
R27
L298
L2
L692
R81
L823
L34
L32
R596
L1
L95
R355
L48
R7
R35
L55
L511
L14
L78
L91
R82
L48
L32
L40
R95
R77
R36
R30
L79
L626
R32
R24
R49
R6
L6
L48
R8
R40
R41
R1
R920
L19
R57
R13
L13
R51
L51
R23
L3
L20
L92
R512
L34
R3
L9
L46
R666
L69
R69
L80
R20
L54
R14
R62
L862
R79
R64
L80
L24
L671
L12
L588
L68
R448
L95
L35
L218
R31
L496
R65
L49
L2
R39
R710
L98
R79
R921
L45
L55
L35
R47
L49
L563
R579
R21
R40
L556
L84
L25
R56
R66
R14
L44
R454
R79
L81
L680
R40
R45
L24
R28
R97
R75
R92
L92
L30
L850
R80
R26
R74
R57
R34
R456
R53
L17
R40
L623
R34
R37
L51
L72
L217
L34
L22
R25
R83
L83
R18
L18
L90
L89
R72
L96
L88
R48
R745
R98
R9
R91
R47
L338
R91
R40
L40
L47
R63
R84
L158
L869
L573
L53
L78
R31
R45
R14
L2
R60
R68
R68
L88
L28
L37
L7
L24
R454
L50
R327
L89
R621
R568
L31
L69
L41
L98
R639
L64
R574
R57
R71
R677
R14
L715
L14
R4
R96
R2
L2
R4
R22
L126
R54
R54
R103
R96
L22
R625
L310
L87
R34
L533
R71
R18
R89
L92
R662
L78
R55
L74
R35
R667
R133
R829
L29
R15
R85
L72
R30
R42
R33
L71
L85
R23
R72
L13
R41
L616
R82
R37
L3
R40
L40
L2
R81
L11
L11
L21
R64
R50
R181
R69
R69
R31
L48
L45
R93
L57
L43
R1
L1
L80
L26
L28
R38
R960
L479
L56
L29
L65
R72
R46
R47
R34
R270
R88
R8
L477
L37
L95
L7
L84
R64
R136
R66
R69
R90
L93
L12
L20
L32
R27
R37
L28
R96
R43
L543
R97
L165
L591
R620
R439
R39
L68
L151
R680
R97
R84
R19
L51
L399
L50
L27
L50
L191
R37
L21
L49
R89
L88
L7
L93
L90
R416
R68
R53
R26
R38
L85
L60
L60
L13
L93
R44
L62
L58
R9
L65
L56
R654
R34
L69
L7
L24
R42
L542
R99
R1
L89
L94
L21
R1
R627
L324
R55
R792
L75
L191
R6
L87
R89
R24
R22
L35
R922
L22
L762
R11
L616
R67
L58
R60
R98
L321
R21
R19
L419
R675
R31
L6
L5
L95
R84
L78
R19
L22
L3
L79
L76
L138
L51
R59
R13
L42
R95
L39
L11
R86
L91
R18
L344
L50
L63
R738
R75
R81
R44
R875
L40
R347
R77
L284
L83
L217
L783
R83
L20
R91
L43
L17
R89
R75
R25
L4
R38
R19
L67
R940
L2
L24
R10
R43
L467
R14
L37
R872
L35
L63
R66
L88
L846
R16
R95
L91
L41
L3
R52
R603
R48
L9
R65
L4
R48
L9
R86
R75
R91
R90
L81
L88
L11
R99
L10
L90
R871
L21
L7
R57
R25
L8
R87
L4
L59
R59
R72
R18
R10
L29
R29
L908
R75
R33
L92
L908
L82
L77
R84
L25
R89
L67
R951
L73
L25
R31
L43
R7
L70
R104
R77
R98
L33
R254
R17
R83
R989
L89
R79
R21
R68
L755
L17
L693
L63
L40
L58
L42
L86
R86
L61
R361
L24
R25
L93
R79
R56
R99
L42
R44
L92
R37
R11
L48
L764
L854
L834
R4
R482
L406
R20
R76
R38
L54
L60
L59
L82
L59
R64
R41
L82
R77
L37
R78
R55
L79
L57
R144
L741
L50
L63
L25
L25
L42
L32
R86
R86
L57
L90
L99
R90
L67
L577
L46
L52
L8
L92
L916
R33
R33
R61
L11
R6
R93
R14
R87
R57
L58
L94
R95
R32
R68
R436
L723
R187
L551
L10
R19
L48
R90
L663
L37
L175
L54
L321
R751
R25
L60
L341
R75
R887
L187
R330
L47
R7
L58
R68
L48
L438
L89
R75
L4
L73
L16
R593
R7
R85
R8
R46
L6
L20
L70
R50
R22
L22
L54
L283
L58
R42
R271
R7
L723
R98
R29
R84
L15
L98
L82
R98
L71
R13
R30
L47
R59
L52
R60
L8
L56
R86
L30
R7
L7
L29
L70
R10
L33
R70
R11
L59
R74
L834
R60
L3
L35
R38
L70
R143
R258
L22
L97
L79
R394
R73
L48
R31
R17
L91
L9
L47
R47
R446
R10
R87
L72
R29
R775
R225
L43
R35
R629
L21
L98
R98
L56
L44
R15
R5
L80
R60
R63
L63
R34
L34
R29
R49
R17
L117
R22
R690
L51
R38
L777
L81
R59
R622
L67
R99
R68
L92
R99
R26
L33
L38
R60
R78
L57
L43
L30
L70
R55
L87
L60
L61
L47
L67
L508
L25
L6
L52
L42
R66
R34
L86
R57
R574
R19
L64
R69
L195
R726
L62
L90
L41
R93
L129
L96
R885
R931
R9
R66
R47
L13
L59
L315
L26
R1
R99
R47
L55
L592
R45
R955
L677
L823
R91
L73
R82
L856
R56
R157
L89
L68
R18
R25
R57
R94
R106
L70
L88
L42
L90
L99
L34
R65
L78
L64
R62
L262
R4
L20
R34
R73
R9
L34
R71
R3
L37
R843
L46
R8
L8
R2
R47
R51
R934
L34
L32
R932
R65
L45
R87
L81
L173
R84
L737
R36
R33
R25
L94
L54
L38
R76
R11
L99
R40
L94
R58
L48
L252
R4
R551
L78
R23
L56
R56
R57
L77
L71
L9
R78
R22
L93
L43
L64
L10
L39
L67
L84
L18
R718
R15
L15
L264
R62
L98
L43
R43
L632
R9
L77
L24
L39
R63
L52
L15
L33
R795
R93
R804
R97
L48
R953
L36
L6
R160
R88
L25
L75
L33
R26
L354
L44
L93
L48
L54
R894
R6
R50
R61
L72
R85
R76
L84
L12
R593
L97
L57
L21
L66
L56
L48
L458
R85
L34
L45
R33
L93
L11
L8
L935
R14
R55
R39
R6
R56
L56
L2
R2
R144
L32
L213
R876
L4
R29
L48
L52
L2
R77
R49
R76
R70
L70
R52
L36
L27
L83
R85
L8
R12
R24
R304
R77
R21
R90
R77
R12
R52
L7
R55
L37
L30
L92
L6
R65
L7
R66
L89
R66
L8
L86
L42
R17
R83
R201
L56
R8
L75
R99
L77
R30
L57
L49
L24
R72
L947
R61
R163
L49
R81
R563
L44
R73
L73
L87
L873
L40
R45
L13
L8
L24
L37
L45
R956
L74
R43
L43
L88
R29
L47
L94
L19
R97
R31
L28
R71
L48
L93
L62
R51
L61
L45
L94
R22
R32
L54
R89
L607
R18
R493
L93
L54
L80
R64
R677
R93
L11
L89
L33
L10
L16
L80
L79
R18
R72
R37
R83
R30
L22
L3
L97
L76
R76
L68
L74
L84
L74
L79
R46
L17
R8
L14
L78
L17
R74
L368
L787
R32
L16
L38
R54
R38
L11
R427
R26
L80
L54
L46
L17
L10
R27
L99
L1
L121
R28
R93
L82
R95
R65
L21
R43
L83
L877
R109
L8
R83
R76
L9
R9
L50
R92
R81
R77
R64
L64
L94
R736
L55
L58
R71
R21
R67
L36
R798
R40
L48
R58
R70
R66
L10
R250
R87
L78
R315
L68
R960
R8
R91
L75
L7
R91
L18
L39
L43
L52
R26
R669
L43
R949
L24
L925
L1
L62
L837
R54
L154
R11
L11
L65
R272
L7
L76
L80
L64
R10
R270
L32
R62
R10
R325
L26
R1
R363
R437
L64
R11
R53
L48
R748
R21
R16
R547
R74
L505
L53
R302
R962
L11
R2
R45
R98
L29
R31
R75
L55
L584
R64
L54
R54
R79
R637
R34
L60
L30
R118
R97
R25
L81
R949
R76
L96
L51
L25
R586
L87
R331
R61
L91
L854
L18
R97
R986
L83
R60
L160
L712
R6
R45
R418
L90
L20
R92
L83
R644
L50
R50
R26
R974
L154
L66
L80
R34
L504
L980
L35
R49
R95
R741
R57
L12
L111
R66
L44
R83
R35
L272
L402
R413
L55
R62
R80
R299
L223
L811
L94
R29
R43
R58
R92
R7
L51
L8
L41
R63
L63
R421
L50
R74
L4
R59
L76
L193
L908
L36
L238
R51
L87
L63
R53
L56
R11
L72
R935
L21
L90
R6
L53
L963
R94
R66
R40
L92
L94
L54
R95
R81
R1
L37
R50
R50
R11
R89
R18
L568
R90
R160
R32
L32
R79
L79
R77
L77
L68
L234
R52
R371
L221
R24
R64
L67
L9
L292
R80
L93
R95
L13
L89
R68
R32
L56
L44
L106
L392
L2
L170
R88
L18
R258
R73
R2
R42
R76
L85
R34
L49
R270
L13
L94
R214
R4
L32
R58
R42
L836
R736
R414
L587
L27
L12
L3
R79
L64
R61
L19
R846
R75
R64
L585
L57
L254
L6
R22
L664
L87
R94
L81
L94
R575
R810
R83
L242
R87
L68
R49
R54
R43
L13
L24
R31
L6
R54
R62
L99
R89
R21
L21
L795
R95
L40
R79
R69
R721
L82
R53
L6
R76
R30
L676
R76
L634
L452
L398
R84
L32
R32
R85
R9
R52
R60
R94
R3
R94
R225
R21
R50
R70
L269
L80
L92
L33
L944
L45
L25
R125
L8
L92
L56
R351
L46
L50
L91
R956
R80
L5
R366
R24
R71
R44
L70
R32
R94
R23
L23
L43
L18
L29
L8
R59
R39
R69
L69
L72
L55
L44
L3
R14
L35
R695
L26
R26
L211
L40
L826
R77
R25
L25
L45
R77
R34
R25
R6
R69
R34
L46
R663
L17
L93
R93
L54
L5
L14
R73
R644
L139
R73
L833
R55
R60
R43
R5
R92
L63
L88
R51
L670
L941
R89
L78
L45
R7
R38
R26
R64
L90
L70
R943
L631
L86
L456
R46
R30
R50
L26
L62
R62
L99
L1
R34
L41
R76
R31
R72
L63
R91
R559
L514
R91
R82
R73
R2
L42
R56
R21
L71
L75
R18
R62
R58
R24
R420
R23
R77
L64
L84
L87
R33
L56
L606
L78
R31
R57
L76
R2
L36
R31
R69
L374
L19
L11
R160
L56
L8
R95
L87
R3
L3
L34
L66
R31
L331
L839
R60
L921
L894
R23
L63
R45
L11
R24
R76
R60
L47
L13
R28
R36
L964
L77
R45
R6
R42
R84
R921
L221
L14
R89
R82
L57
R65
L591
L725
L49
L922
R22
R64
R307
L96
R13
R12
R84
L212
L772
L7
L346
R46
L46
R45
L592
R80
R145
L93
L214
R82
L696
L4
L58
R30
R89
R45
L34
L72
R86
L38
L48
L35
R7
R28
R63
L63
R46
L46
R38
L38
R12
R93
L47
R42
L55
R23
R77
R55
R56
R547
L86
R83
R87
R73
R50
R35
R55
R54
L89
R88
R57
R90
L19
R43
L24
L70
L30
L1
L97
R81
L95
R81
R16
L85
L89
R60
R7
L47
R69
R45
L45
L97
R97
L47
L53
L12
L1
R13
R37
R87
R67
L54
R63
R96
R4
R65
R63
L28
R70
L20
L55
R72
R59
R62
L78
R89
L87
R88
R54
R46
R70
L70
R63
L63
R12
L12
L99
R99
R46
L46
L36
R7
L12
L5
L31
L34
R36
R42
R41
L10
R17
L21
R18
L16
L33
L9
L33
L13
L50
L36
R20
R15
L29
R16
R31
L2
L12
L40
R41
R47
R8
L42
L48
R45
L29
R42
R20
L33
L7
R22
R32
L20
L14
L28
L17
R33
R6
R39
R47
R9
L5";
        
        // Temporary variables for parsing
        byte dir_char0, dir_char1;  // For 'R' or 'L'
        integer mag0, mag1;         // For numbers
        integer scan_result;
        
        // Parse the string using $sscanf
        scan_result = $sscanf(input_str, "%c%d %c%d", dir_char0, mag0, dir_char1, mag1);
        
        // Check if parsing succeeded (should match 4 items)
        if (scan_result != 4) begin
            $display("Error: Parsing failed! Check input string format.");
            $finish;
        end
        
        // Map characters to 0/1
        direction[0] = (dir_char0 == "R") ? 1'b0 : 1'b1;
        direction[1] = (dir_char1 == "L") ? 1'b1 : 1'b0;
        
        // Assign magnitudes directly
        magnitude[0] = mag0;
        magnitude[1] = mag1;
        
        // Display the results
        $display("Direction vector: [%0d, %0d]", direction[0], direction[1]);
        $display("Magnitude vector: [%0d, %0d]", magnitude[0], magnitude[1]);
        
        // End simulation
        $finish;
    end

endmodule